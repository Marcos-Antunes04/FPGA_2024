NET "BUT[0]" CLOCK_DEDICATED_ROUTE = FALSE;

NET "CLK27MHz" LOC = V10 ;

NET "GPIO[0]" LOC = N17;
NET "GPIO[1]" LOC = M18;
NET "GPIO[2]" LOC = A3;
NET "GPIO[3]" LOC = L15;
NET "GPIO[4]" LOC = F15;
NET "GPIO[5]" LOC = B4;
NET "GPIO[6]" LOC = F13;
NET "GPIO[7]" LOC = P12;

NET "BUT[0]" LOC = P4;
NET "BUT[1]" LOC = F6;
NET "BUT[2]" LOC = E4;
NET "BUT[3]" LOC = F5;

NET "DIPSW[0]" LOC = D14;
NET "DIPSW[1]" LOC = E12;
NET "DIPSW[2]" LOC = F12;
NET "DIPSW[3]" LOC = V13;

NET "LEDS[0]" LOC = E13;
NET "LEDS[1]" LOC = C14;
NET "LEDS[2]" LOC = C4;
NET "LEDS[3]" LOC = A4;