library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity flip-flop-D is port ();
end flip-flop-D;

architecture Hardware of flip-flop-D is

begin


end Hardware;

